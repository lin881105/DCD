module Lab2_BCD_3bit_add(BCD_X,BCD_Y,cin,BCD_S,cout);
input   [11:0]   BCD_X,BCD_Y;
output  [11:0]   BCD_S;
input           cin;
output          cout;
wire            cout1,cout2;

Lab2_BCD_1bit_add_beh		M1(BCD_X[3:0], BCD_Y[3:0], cin,BCD_S[3:0],cout1);
Lab2_BCD_1bit_add_beh		M2(BCD_X[7:4], BCD_Y[7:4], cout1,BCD_S[7:4],cout2);
Lab2_BCD_1bit_add_beh		M3(BCD_X[11:8], BCD_Y[11:8], cout2,BCD_S[11:8],cout);

endmodule